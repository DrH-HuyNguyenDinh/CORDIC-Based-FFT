module rom_stage_9 (
    input logic         i_clk,
    input logic [7:0]   i_addr,   
    output logic [31:0] o_data
);

logic [31:0] rom [0:255];

initial begin
    rom[  0] = 32'h80000000; // 0 * -pi/256 (-0.00 deg)
    rom[  1] = 32'hbc490fdb; // 1 * -pi/256 (-0.70 deg)
    rom[  2] = 32'hbcc90fdb; // 2 * -pi/256 (-1.41 deg)
    rom[  3] = 32'hbd16cbe4; // 3 * -pi/256 (-2.11 deg)
    rom[  4] = 32'hbd490fdb; // 4 * -pi/256 (-2.81 deg)
    rom[  5] = 32'hbd7b53d1; // 5 * -pi/256 (-3.52 deg)
    rom[  6] = 32'hbd96cbe4; // 6 * -pi/256 (-4.22 deg)
    rom[  7] = 32'hbdafeddf; // 7 * -pi/256 (-4.92 deg)
    rom[  8] = 32'hbdc90fdb; // 8 * -pi/256 (-5.62 deg)
    rom[  9] = 32'hbde231d6; // 9 * -pi/256 (-6.33 deg)
    rom[ 10] = 32'hbdfb53d1; // 10 * -pi/256 (-7.03 deg)
    rom[ 11] = 32'hbe0a3ae6; // 11 * -pi/256 (-7.73 deg)
    rom[ 12] = 32'hbe16cbe4; // 12 * -pi/256 (-8.44 deg)
    rom[ 13] = 32'hbe235ce2; // 13 * -pi/256 (-9.14 deg)
    rom[ 14] = 32'hbe2feddf; // 14 * -pi/256 (-9.84 deg)
    rom[ 15] = 32'hbe3c7edd; // 15 * -pi/256 (-10.55 deg)
    rom[ 16] = 32'hbe490fdb; // 16 * -pi/256 (-11.25 deg)
    rom[ 17] = 32'hbe55a0d8; // 17 * -pi/256 (-11.95 deg)
    rom[ 18] = 32'hbe6231d6; // 18 * -pi/256 (-12.66 deg)
    rom[ 19] = 32'hbe6ec2d4; // 19 * -pi/256 (-13.36 deg)
    rom[ 20] = 32'hbe7b53d1; // 20 * -pi/256 (-14.06 deg)
    rom[ 21] = 32'hbe83f267; // 21 * -pi/256 (-14.77 deg)
    rom[ 22] = 32'hbe8a3ae6; // 22 * -pi/256 (-15.47 deg)
    rom[ 23] = 32'hbe908365; // 23 * -pi/256 (-16.17 deg)
    rom[ 24] = 32'hbe96cbe4; // 24 * -pi/256 (-16.88 deg)
    rom[ 25] = 32'hbe9d1463; // 25 * -pi/256 (-17.58 deg)
    rom[ 26] = 32'hbea35ce2; // 26 * -pi/256 (-18.28 deg)
    rom[ 27] = 32'hbea9a560; // 27 * -pi/256 (-18.98 deg)
    rom[ 28] = 32'hbeafeddf; // 28 * -pi/256 (-19.69 deg)
    rom[ 29] = 32'hbeb6365e; // 29 * -pi/256 (-20.39 deg)
    rom[ 30] = 32'hbebc7edd; // 30 * -pi/256 (-21.09 deg)
    rom[ 31] = 32'hbec2c75c; // 31 * -pi/256 (-21.80 deg)
    rom[ 32] = 32'hbec90fdb; // 32 * -pi/256 (-22.50 deg)
    rom[ 33] = 32'hbecf5859; // 33 * -pi/256 (-23.20 deg)
    rom[ 34] = 32'hbed5a0d8; // 34 * -pi/256 (-23.91 deg)
    rom[ 35] = 32'hbedbe957; // 35 * -pi/256 (-24.61 deg)
    rom[ 36] = 32'hbee231d6; // 36 * -pi/256 (-25.31 deg)
    rom[ 37] = 32'hbee87a55; // 37 * -pi/256 (-26.02 deg)
    rom[ 38] = 32'hbeeec2d4; // 38 * -pi/256 (-26.72 deg)
    rom[ 39] = 32'hbef50b52; // 39 * -pi/256 (-27.42 deg)
    rom[ 40] = 32'hbefb53d1; // 40 * -pi/256 (-28.12 deg)
    rom[ 41] = 32'hbf00ce28; // 41 * -pi/256 (-28.83 deg)
    rom[ 42] = 32'hbf03f267; // 42 * -pi/256 (-29.53 deg)
    rom[ 43] = 32'hbf0716a7; // 43 * -pi/256 (-30.23 deg)
    rom[ 44] = 32'hbf0a3ae6; // 44 * -pi/256 (-30.94 deg)
    rom[ 45] = 32'hbf0d5f26; // 45 * -pi/256 (-31.64 deg)
    rom[ 46] = 32'hbf108365; // 46 * -pi/256 (-32.34 deg)
    rom[ 47] = 32'hbf13a7a5; // 47 * -pi/256 (-33.05 deg)
    rom[ 48] = 32'hbf16cbe4; // 48 * -pi/256 (-33.75 deg)
    rom[ 49] = 32'hbf19f023; // 49 * -pi/256 (-34.45 deg)
    rom[ 50] = 32'hbf1d1463; // 50 * -pi/256 (-35.16 deg)
    rom[ 51] = 32'hbf2038a2; // 51 * -pi/256 (-35.86 deg)
    rom[ 52] = 32'hbf235ce2; // 52 * -pi/256 (-36.56 deg)
    rom[ 53] = 32'hbf268121; // 53 * -pi/256 (-37.27 deg)
    rom[ 54] = 32'hbf29a560; // 54 * -pi/256 (-37.97 deg)
    rom[ 55] = 32'hbf2cc9a0; // 55 * -pi/256 (-38.67 deg)
    rom[ 56] = 32'hbf2feddf; // 56 * -pi/256 (-39.38 deg)
    rom[ 57] = 32'hbf33121f; // 57 * -pi/256 (-40.08 deg)
    rom[ 58] = 32'hbf36365e; // 58 * -pi/256 (-40.78 deg)
    rom[ 59] = 32'hbf395a9e; // 59 * -pi/256 (-41.48 deg)
    rom[ 60] = 32'hbf3c7edd; // 60 * -pi/256 (-42.19 deg)
    rom[ 61] = 32'hbf3fa31c; // 61 * -pi/256 (-42.89 deg)
    rom[ 62] = 32'hbf42c75c; // 62 * -pi/256 (-43.59 deg)
    rom[ 63] = 32'hbf45eb9b; // 63 * -pi/256 (-44.30 deg)
    rom[ 64] = 32'hbf490fdb; // 64 * -pi/256 (-45.00 deg)
    rom[ 65] = 32'hbf4c341a; // 65 * -pi/256 (-45.70 deg)
    rom[ 66] = 32'hbf4f5859; // 66 * -pi/256 (-46.41 deg)
    rom[ 67] = 32'hbf527c99; // 67 * -pi/256 (-47.11 deg)
    rom[ 68] = 32'hbf55a0d8; // 68 * -pi/256 (-47.81 deg)
    rom[ 69] = 32'hbf58c518; // 69 * -pi/256 (-48.52 deg)
    rom[ 70] = 32'hbf5be957; // 70 * -pi/256 (-49.22 deg)
    rom[ 71] = 32'hbf5f0d97; // 71 * -pi/256 (-49.92 deg)
    rom[ 72] = 32'hbf6231d6; // 72 * -pi/256 (-50.62 deg)
    rom[ 73] = 32'hbf655615; // 73 * -pi/256 (-51.33 deg)
    rom[ 74] = 32'hbf687a55; // 74 * -pi/256 (-52.03 deg)
    rom[ 75] = 32'hbf6b9e94; // 75 * -pi/256 (-52.73 deg)
    rom[ 76] = 32'hbf6ec2d4; // 76 * -pi/256 (-53.44 deg)
    rom[ 77] = 32'hbf71e713; // 77 * -pi/256 (-54.14 deg)
    rom[ 78] = 32'hbf750b52; // 78 * -pi/256 (-54.84 deg)
    rom[ 79] = 32'hbf782f92; // 79 * -pi/256 (-55.55 deg)
    rom[ 80] = 32'hbf7b53d1; // 80 * -pi/256 (-56.25 deg)
    rom[ 81] = 32'hbf7e7811; // 81 * -pi/256 (-56.95 deg)
    rom[ 82] = 32'hbf80ce28; // 82 * -pi/256 (-57.66 deg)
    rom[ 83] = 32'hbf826048; // 83 * -pi/256 (-58.36 deg)
    rom[ 84] = 32'hbf83f267; // 84 * -pi/256 (-59.06 deg)
    rom[ 85] = 32'hbf858487; // 85 * -pi/256 (-59.77 deg)
    rom[ 86] = 32'hbf8716a7; // 86 * -pi/256 (-60.47 deg)
    rom[ 87] = 32'hbf88a8c7; // 87 * -pi/256 (-61.17 deg)
    rom[ 88] = 32'hbf8a3ae6; // 88 * -pi/256 (-61.87 deg)
    rom[ 89] = 32'hbf8bcd06; // 89 * -pi/256 (-62.58 deg)
    rom[ 90] = 32'hbf8d5f26; // 90 * -pi/256 (-63.28 deg)
    rom[ 91] = 32'hbf8ef145; // 91 * -pi/256 (-63.98 deg)
    rom[ 92] = 32'hbf908365; // 92 * -pi/256 (-64.69 deg)
    rom[ 93] = 32'hbf921585; // 93 * -pi/256 (-65.39 deg)
    rom[ 94] = 32'hbf93a7a5; // 94 * -pi/256 (-66.09 deg)
    rom[ 95] = 32'hbf9539c4; // 95 * -pi/256 (-66.80 deg)
    rom[ 96] = 32'hbf96cbe4; // 96 * -pi/256 (-67.50 deg)
    rom[ 97] = 32'hbf985e04; // 97 * -pi/256 (-68.20 deg)
    rom[ 98] = 32'hbf99f023; // 98 * -pi/256 (-68.91 deg)
    rom[ 99] = 32'hbf9b8243; // 99 * -pi/256 (-69.61 deg)
    rom[100] = 32'hbf9d1463; // 100 * -pi/256 (-70.31 deg)
    rom[101] = 32'hbf9ea683; // 101 * -pi/256 (-71.02 deg)
    rom[102] = 32'hbfa038a2; // 102 * -pi/256 (-71.72 deg)
    rom[103] = 32'hbfa1cac2; // 103 * -pi/256 (-72.42 deg)
    rom[104] = 32'hbfa35ce2; // 104 * -pi/256 (-73.12 deg)
    rom[105] = 32'hbfa4ef01; // 105 * -pi/256 (-73.83 deg)
    rom[106] = 32'hbfa68121; // 106 * -pi/256 (-74.53 deg)
    rom[107] = 32'hbfa81341; // 107 * -pi/256 (-75.23 deg)
    rom[108] = 32'hbfa9a560; // 108 * -pi/256 (-75.94 deg)
    rom[109] = 32'hbfab3780; // 109 * -pi/256 (-76.64 deg)
    rom[110] = 32'hbfacc9a0; // 110 * -pi/256 (-77.34 deg)
    rom[111] = 32'hbfae5bc0; // 111 * -pi/256 (-78.05 deg)
    rom[112] = 32'hbfafeddf; // 112 * -pi/256 (-78.75 deg)
    rom[113] = 32'hbfb17fff; // 113 * -pi/256 (-79.45 deg)
    rom[114] = 32'hbfb3121f; // 114 * -pi/256 (-80.16 deg)
    rom[115] = 32'hbfb4a43e; // 115 * -pi/256 (-80.86 deg)
    rom[116] = 32'hbfb6365e; // 116 * -pi/256 (-81.56 deg)
    rom[117] = 32'hbfb7c87e; // 117 * -pi/256 (-82.27 deg)
    rom[118] = 32'hbfb95a9e; // 118 * -pi/256 (-82.97 deg)
    rom[119] = 32'hbfbaecbd; // 119 * -pi/256 (-83.67 deg)
    rom[120] = 32'hbfbc7edd; // 120 * -pi/256 (-84.38 deg)
    rom[121] = 32'hbfbe10fd; // 121 * -pi/256 (-85.08 deg)
    rom[122] = 32'hbfbfa31c; // 122 * -pi/256 (-85.78 deg)
    rom[123] = 32'hbfc1353c; // 123 * -pi/256 (-86.48 deg)
    rom[124] = 32'hbfc2c75c; // 124 * -pi/256 (-87.19 deg)
    rom[125] = 32'hbfc4597c; // 125 * -pi/256 (-87.89 deg)
    rom[126] = 32'hbfc5eb9b; // 126 * -pi/256 (-88.59 deg)
    rom[127] = 32'hbfc77dbb; // 127 * -pi/256 (-89.30 deg)
    rom[128] = 32'hbfc90fdb; // 128 * -pi/256 (-90.00 deg)
    rom[129] = 32'hbfcaa1fa; // 129 * -pi/256 (-90.70 deg)
    rom[130] = 32'hbfcc341a; // 130 * -pi/256 (-91.41 deg)
    rom[131] = 32'hbfcdc63a; // 131 * -pi/256 (-92.11 deg)
    rom[132] = 32'hbfcf5859; // 132 * -pi/256 (-92.81 deg)
    rom[133] = 32'hbfd0ea79; // 133 * -pi/256 (-93.52 deg)
    rom[134] = 32'hbfd27c99; // 134 * -pi/256 (-94.22 deg)
    rom[135] = 32'hbfd40eb9; // 135 * -pi/256 (-94.92 deg)
    rom[136] = 32'hbfd5a0d8; // 136 * -pi/256 (-95.62 deg)
    rom[137] = 32'hbfd732f8; // 137 * -pi/256 (-96.33 deg)
    rom[138] = 32'hbfd8c518; // 138 * -pi/256 (-97.03 deg)
    rom[139] = 32'hbfda5737; // 139 * -pi/256 (-97.73 deg)
    rom[140] = 32'hbfdbe957; // 140 * -pi/256 (-98.44 deg)
    rom[141] = 32'hbfdd7b77; // 141 * -pi/256 (-99.14 deg)
    rom[142] = 32'hbfdf0d97; // 142 * -pi/256 (-99.84 deg)
    rom[143] = 32'hbfe09fb6; // 143 * -pi/256 (-100.55 deg)
    rom[144] = 32'hbfe231d6; // 144 * -pi/256 (-101.25 deg)
    rom[145] = 32'hbfe3c3f6; // 145 * -pi/256 (-101.95 deg)
    rom[146] = 32'hbfe55615; // 146 * -pi/256 (-102.66 deg)
    rom[147] = 32'hbfe6e835; // 147 * -pi/256 (-103.36 deg)
    rom[148] = 32'hbfe87a55; // 148 * -pi/256 (-104.06 deg)
    rom[149] = 32'hbfea0c75; // 149 * -pi/256 (-104.77 deg)
    rom[150] = 32'hbfeb9e94; // 150 * -pi/256 (-105.47 deg)
    rom[151] = 32'hbfed30b4; // 151 * -pi/256 (-106.17 deg)
    rom[152] = 32'hbfeec2d4; // 152 * -pi/256 (-106.88 deg)
    rom[153] = 32'hbff054f3; // 153 * -pi/256 (-107.58 deg)
    rom[154] = 32'hbff1e713; // 154 * -pi/256 (-108.28 deg)
    rom[155] = 32'hbff37933; // 155 * -pi/256 (-108.98 deg)
    rom[156] = 32'hbff50b52; // 156 * -pi/256 (-109.69 deg)
    rom[157] = 32'hbff69d72; // 157 * -pi/256 (-110.39 deg)
    rom[158] = 32'hbff82f92; // 158 * -pi/256 (-111.09 deg)
    rom[159] = 32'hbff9c1b2; // 159 * -pi/256 (-111.80 deg)
    rom[160] = 32'hbffb53d1; // 160 * -pi/256 (-112.50 deg)
    rom[161] = 32'hbffce5f1; // 161 * -pi/256 (-113.20 deg)
    rom[162] = 32'hbffe7811; // 162 * -pi/256 (-113.91 deg)
    rom[163] = 32'hc0000518; // 163 * -pi/256 (-114.61 deg)
    rom[164] = 32'hc000ce28; // 164 * -pi/256 (-115.31 deg)
    rom[165] = 32'hc0019738; // 165 * -pi/256 (-116.02 deg)
    rom[166] = 32'hc0026048; // 166 * -pi/256 (-116.72 deg)
    rom[167] = 32'hc0032958; // 167 * -pi/256 (-117.42 deg)
    rom[168] = 32'hc003f267; // 168 * -pi/256 (-118.12 deg)
    rom[169] = 32'hc004bb77; // 169 * -pi/256 (-118.83 deg)
    rom[170] = 32'hc0058487; // 170 * -pi/256 (-119.53 deg)
    rom[171] = 32'hc0064d97; // 171 * -pi/256 (-120.23 deg)
    rom[172] = 32'hc00716a7; // 172 * -pi/256 (-120.94 deg)
    rom[173] = 32'hc007dfb7; // 173 * -pi/256 (-121.64 deg)
    rom[174] = 32'hc008a8c7; // 174 * -pi/256 (-122.34 deg)
    rom[175] = 32'hc00971d6; // 175 * -pi/256 (-123.05 deg)
    rom[176] = 32'hc00a3ae6; // 176 * -pi/256 (-123.75 deg)
    rom[177] = 32'hc00b03f6; // 177 * -pi/256 (-124.45 deg)
    rom[178] = 32'hc00bcd06; // 178 * -pi/256 (-125.16 deg)
    rom[179] = 32'hc00c9616; // 179 * -pi/256 (-125.86 deg)
    rom[180] = 32'hc00d5f26; // 180 * -pi/256 (-126.56 deg)
    rom[181] = 32'hc00e2836; // 181 * -pi/256 (-127.27 deg)
    rom[182] = 32'hc00ef145; // 182 * -pi/256 (-127.97 deg)
    rom[183] = 32'hc00fba55; // 183 * -pi/256 (-128.67 deg)
    rom[184] = 32'hc0108365; // 184 * -pi/256 (-129.38 deg)
    rom[185] = 32'hc0114c75; // 185 * -pi/256 (-130.08 deg)
    rom[186] = 32'hc0121585; // 186 * -pi/256 (-130.78 deg)
    rom[187] = 32'hc012de95; // 187 * -pi/256 (-131.48 deg)
    rom[188] = 32'hc013a7a5; // 188 * -pi/256 (-132.19 deg)
    rom[189] = 32'hc01470b4; // 189 * -pi/256 (-132.89 deg)
    rom[190] = 32'hc01539c4; // 190 * -pi/256 (-133.59 deg)
    rom[191] = 32'hc01602d4; // 191 * -pi/256 (-134.30 deg)
    rom[192] = 32'hc016cbe4; // 192 * -pi/256 (-135.00 deg)
    rom[193] = 32'hc01794f4; // 193 * -pi/256 (-135.70 deg)
    rom[194] = 32'hc0185e04; // 194 * -pi/256 (-136.41 deg)
    rom[195] = 32'hc0192714; // 195 * -pi/256 (-137.11 deg)
    rom[196] = 32'hc019f023; // 196 * -pi/256 (-137.81 deg)
    rom[197] = 32'hc01ab933; // 197 * -pi/256 (-138.52 deg)
    rom[198] = 32'hc01b8243; // 198 * -pi/256 (-139.22 deg)
    rom[199] = 32'hc01c4b53; // 199 * -pi/256 (-139.92 deg)
    rom[200] = 32'hc01d1463; // 200 * -pi/256 (-140.62 deg)
    rom[201] = 32'hc01ddd73; // 201 * -pi/256 (-141.33 deg)
    rom[202] = 32'hc01ea683; // 202 * -pi/256 (-142.03 deg)
    rom[203] = 32'hc01f6f92; // 203 * -pi/256 (-142.73 deg)
    rom[204] = 32'hc02038a2; // 204 * -pi/256 (-143.44 deg)
    rom[205] = 32'hc02101b2; // 205 * -pi/256 (-144.14 deg)
    rom[206] = 32'hc021cac2; // 206 * -pi/256 (-144.84 deg)
    rom[207] = 32'hc02293d2; // 207 * -pi/256 (-145.55 deg)
    rom[208] = 32'hc0235ce2; // 208 * -pi/256 (-146.25 deg)
    rom[209] = 32'hc02425f1; // 209 * -pi/256 (-146.95 deg)
    rom[210] = 32'hc024ef01; // 210 * -pi/256 (-147.66 deg)
    rom[211] = 32'hc025b811; // 211 * -pi/256 (-148.36 deg)
    rom[212] = 32'hc0268121; // 212 * -pi/256 (-149.06 deg)
    rom[213] = 32'hc0274a31; // 213 * -pi/256 (-149.77 deg)
    rom[214] = 32'hc0281341; // 214 * -pi/256 (-150.47 deg)
    rom[215] = 32'hc028dc51; // 215 * -pi/256 (-151.17 deg)
    rom[216] = 32'hc029a560; // 216 * -pi/256 (-151.88 deg)
    rom[217] = 32'hc02a6e70; // 217 * -pi/256 (-152.58 deg)
    rom[218] = 32'hc02b3780; // 218 * -pi/256 (-153.28 deg)
    rom[219] = 32'hc02c0090; // 219 * -pi/256 (-153.98 deg)
    rom[220] = 32'hc02cc9a0; // 220 * -pi/256 (-154.69 deg)
    rom[221] = 32'hc02d92b0; // 221 * -pi/256 (-155.39 deg)
    rom[222] = 32'hc02e5bc0; // 222 * -pi/256 (-156.09 deg)
    rom[223] = 32'hc02f24cf; // 223 * -pi/256 (-156.80 deg)
    rom[224] = 32'hc02feddf; // 224 * -pi/256 (-157.50 deg)
    rom[225] = 32'hc030b6ef; // 225 * -pi/256 (-158.20 deg)
    rom[226] = 32'hc0317fff; // 226 * -pi/256 (-158.91 deg)
    rom[227] = 32'hc032490f; // 227 * -pi/256 (-159.61 deg)
    rom[228] = 32'hc033121f; // 228 * -pi/256 (-160.31 deg)
    rom[229] = 32'hc033db2f; // 229 * -pi/256 (-161.02 deg)
    rom[230] = 32'hc034a43e; // 230 * -pi/256 (-161.72 deg)
    rom[231] = 32'hc0356d4e; // 231 * -pi/256 (-162.42 deg)
    rom[232] = 32'hc036365e; // 232 * -pi/256 (-163.12 deg)
    rom[233] = 32'hc036ff6e; // 233 * -pi/256 (-163.83 deg)
    rom[234] = 32'hc037c87e; // 234 * -pi/256 (-164.53 deg)
    rom[235] = 32'hc038918e; // 235 * -pi/256 (-165.23 deg)
    rom[236] = 32'hc0395a9e; // 236 * -pi/256 (-165.94 deg)
    rom[237] = 32'hc03a23ad; // 237 * -pi/256 (-166.64 deg)
    rom[238] = 32'hc03aecbd; // 238 * -pi/256 (-167.34 deg)
    rom[239] = 32'hc03bb5cd; // 239 * -pi/256 (-168.05 deg)
    rom[240] = 32'hc03c7edd; // 240 * -pi/256 (-168.75 deg)
    rom[241] = 32'hc03d47ed; // 241 * -pi/256 (-169.45 deg)
    rom[242] = 32'hc03e10fd; // 242 * -pi/256 (-170.16 deg)
    rom[243] = 32'hc03eda0d; // 243 * -pi/256 (-170.86 deg)
    rom[244] = 32'hc03fa31c; // 244 * -pi/256 (-171.56 deg)
    rom[245] = 32'hc0406c2c; // 245 * -pi/256 (-172.27 deg)
    rom[246] = 32'hc041353c; // 246 * -pi/256 (-172.97 deg)
    rom[247] = 32'hc041fe4c; // 247 * -pi/256 (-173.67 deg)
    rom[248] = 32'hc042c75c; // 248 * -pi/256 (-174.38 deg)
    rom[249] = 32'hc043906c; // 249 * -pi/256 (-175.08 deg)
    rom[250] = 32'hc044597c; // 250 * -pi/256 (-175.78 deg)
    rom[251] = 32'hc045228b; // 251 * -pi/256 (-176.48 deg)
    rom[252] = 32'hc045eb9b; // 252 * -pi/256 (-177.19 deg)
    rom[253] = 32'hc046b4ab; // 253 * -pi/256 (-177.89 deg)
    rom[254] = 32'hc0477dbb; // 254 * -pi/256 (-178.59 deg)
    rom[255] = 32'hc04846cb; // 255 * -pi/256 (-179.30 deg)
end

always @(posedge i_clk) begin
    o_data <= rom[i_addr];
end

endmodule
