module rom_stage_10 (
    input logic         i_clk,
    input logic [8:0]   i_addr,   // [THAY ĐỔI]: 9 bit cho 512 góc
    output logic [31:0] o_data
);

logic [31:0] rom [0:511];

initial begin
    rom[  0] = 32'h80000000; // 0 * -pi/512
    rom[  1] = 32'hbbc90fdb; // 1 * -pi/512
    rom[  2] = 32'hbc490fdb; // 2 * -pi/512
    rom[  3] = 32'hbc96cbe4; // 3 * -pi/512
    rom[  4] = 32'hbcc90fdb; // 4 * -pi/512
    rom[  5] = 32'hbcfb53d1; // 5 * -pi/512
    rom[  6] = 32'hbd16cbe4; // 6 * -pi/512
    rom[  7] = 32'hbd2feddf; // 7 * -pi/512
    rom[  8] = 32'hbd490fdb; // 8 * -pi/512
    rom[  9] = 32'hbd6231d6; // 9 * -pi/512
    rom[ 10] = 32'hbd7b53d1; // 10 * -pi/512
    rom[ 11] = 32'hbd8a3ae6; // 11 * -pi/512
    rom[ 12] = 32'hbd96cbe4; // 12 * -pi/512
    rom[ 13] = 32'hbda35ce2; // 13 * -pi/512
    rom[ 14] = 32'hbdafeddf; // 14 * -pi/512
    rom[ 15] = 32'hbdbc7edd; // 15 * -pi/512
    rom[ 16] = 32'hbdc90fdb; // 16 * -pi/512
    rom[ 17] = 32'hbdd5a0d8; // 17 * -pi/512
    rom[ 18] = 32'hbde231d6; // 18 * -pi/512
    rom[ 19] = 32'hbdeec2d4; // 19 * -pi/512
    rom[ 20] = 32'hbdfb53d1; // 20 * -pi/512
    rom[ 21] = 32'hbe03f267; // 21 * -pi/512
    rom[ 22] = 32'hbe0a3ae6; // 22 * -pi/512
    rom[ 23] = 32'hbe108365; // 23 * -pi/512
    rom[ 24] = 32'hbe16cbe4; // 24 * -pi/512
    rom[ 25] = 32'hbe1d1463; // 25 * -pi/512
    rom[ 26] = 32'hbe235ce2; // 26 * -pi/512
    rom[ 27] = 32'hbe29a560; // 27 * -pi/512
    rom[ 28] = 32'hbe2feddf; // 28 * -pi/512
    rom[ 29] = 32'hbe36365e; // 29 * -pi/512
    rom[ 30] = 32'hbe3c7edd; // 30 * -pi/512
    rom[ 31] = 32'hbe42c75c; // 31 * -pi/512
    rom[ 32] = 32'hbe490fdb; // 32 * -pi/512
    rom[ 33] = 32'hbe4f5859; // 33 * -pi/512
    rom[ 34] = 32'hbe55a0d8; // 34 * -pi/512
    rom[ 35] = 32'hbe5be957; // 35 * -pi/512
    rom[ 36] = 32'hbe6231d6; // 36 * -pi/512
    rom[ 37] = 32'hbe687a55; // 37 * -pi/512
    rom[ 38] = 32'hbe6ec2d4; // 38 * -pi/512
    rom[ 39] = 32'hbe750b52; // 39 * -pi/512
    rom[ 40] = 32'hbe7b53d1; // 40 * -pi/512
    rom[ 41] = 32'hbe80ce28; // 41 * -pi/512
    rom[ 42] = 32'hbe83f267; // 42 * -pi/512
    rom[ 43] = 32'hbe8716a7; // 43 * -pi/512
    rom[ 44] = 32'hbe8a3ae6; // 44 * -pi/512
    rom[ 45] = 32'hbe8d5f26; // 45 * -pi/512
    rom[ 46] = 32'hbe908365; // 46 * -pi/512
    rom[ 47] = 32'hbe93a7a5; // 47 * -pi/512
    rom[ 48] = 32'hbe96cbe4; // 48 * -pi/512
    rom[ 49] = 32'hbe99f023; // 49 * -pi/512
    rom[ 50] = 32'hbe9d1463; // 50 * -pi/512
    rom[ 51] = 32'hbea038a2; // 51 * -pi/512
    rom[ 52] = 32'hbea35ce2; // 52 * -pi/512
    rom[ 53] = 32'hbea68121; // 53 * -pi/512
    rom[ 54] = 32'hbea9a560; // 54 * -pi/512
    rom[ 55] = 32'hbeacc9a0; // 55 * -pi/512
    rom[ 56] = 32'hbeafeddf; // 56 * -pi/512
    rom[ 57] = 32'hbeb3121f; // 57 * -pi/512
    rom[ 58] = 32'hbeb6365e; // 58 * -pi/512
    rom[ 59] = 32'hbeb95a9e; // 59 * -pi/512
    rom[ 60] = 32'hbebc7edd; // 60 * -pi/512
    rom[ 61] = 32'hbebfa31c; // 61 * -pi/512
    rom[ 62] = 32'hbec2c75c; // 62 * -pi/512
    rom[ 63] = 32'hbec5eb9b; // 63 * -pi/512
    rom[ 64] = 32'hbec90fdb; // 64 * -pi/512
    rom[ 65] = 32'hbecc341a; // 65 * -pi/512
    rom[ 66] = 32'hbecf5859; // 66 * -pi/512
    rom[ 67] = 32'hbed27c99; // 67 * -pi/512
    rom[ 68] = 32'hbed5a0d8; // 68 * -pi/512
    rom[ 69] = 32'hbed8c518; // 69 * -pi/512
    rom[ 70] = 32'hbedbe957; // 70 * -pi/512
    rom[ 71] = 32'hbedf0d97; // 71 * -pi/512
    rom[ 72] = 32'hbee231d6; // 72 * -pi/512
    rom[ 73] = 32'hbee55615; // 73 * -pi/512
    rom[ 74] = 32'hbee87a55; // 74 * -pi/512
    rom[ 75] = 32'hbeeb9e94; // 75 * -pi/512
    rom[ 76] = 32'hbeeec2d4; // 76 * -pi/512
    rom[ 77] = 32'hbef1e713; // 77 * -pi/512
    rom[ 78] = 32'hbef50b52; // 78 * -pi/512
    rom[ 79] = 32'hbef82f92; // 79 * -pi/512
    rom[ 80] = 32'hbefb53d1; // 80 * -pi/512
    rom[ 81] = 32'hbefe7811; // 81 * -pi/512
    rom[ 82] = 32'hbf00ce28; // 82 * -pi/512
    rom[ 83] = 32'hbf026048; // 83 * -pi/512
    rom[ 84] = 32'hbf03f267; // 84 * -pi/512
    rom[ 85] = 32'hbf058487; // 85 * -pi/512
    rom[ 86] = 32'hbf0716a7; // 86 * -pi/512
    rom[ 87] = 32'hbf08a8c7; // 87 * -pi/512
    rom[ 88] = 32'hbf0a3ae6; // 88 * -pi/512
    rom[ 89] = 32'hbf0bcd06; // 89 * -pi/512
    rom[ 90] = 32'hbf0d5f26; // 90 * -pi/512
    rom[ 91] = 32'hbf0ef145; // 91 * -pi/512
    rom[ 92] = 32'hbf108365; // 92 * -pi/512
    rom[ 93] = 32'hbf121585; // 93 * -pi/512
    rom[ 94] = 32'hbf13a7a5; // 94 * -pi/512
    rom[ 95] = 32'hbf1539c4; // 95 * -pi/512
    rom[ 96] = 32'hbf16cbe4; // 96 * -pi/512
    rom[ 97] = 32'hbf185e04; // 97 * -pi/512
    rom[ 98] = 32'hbf19f023; // 98 * -pi/512
    rom[ 99] = 32'hbf1b8243; // 99 * -pi/512
    rom[100] = 32'hbf1d1463; // 100 * -pi/512
    rom[101] = 32'hbf1ea683; // 101 * -pi/512
    rom[102] = 32'hbf2038a2; // 102 * -pi/512
    rom[103] = 32'hbf21cac2; // 103 * -pi/512
    rom[104] = 32'hbf235ce2; // 104 * -pi/512
    rom[105] = 32'hbf24ef01; // 105 * -pi/512
    rom[106] = 32'hbf268121; // 106 * -pi/512
    rom[107] = 32'hbf281341; // 107 * -pi/512
    rom[108] = 32'hbf29a560; // 108 * -pi/512
    rom[109] = 32'hbf2b3780; // 109 * -pi/512
    rom[110] = 32'hbf2cc9a0; // 110 * -pi/512
    rom[111] = 32'hbf2e5bc0; // 111 * -pi/512
    rom[112] = 32'hbf2feddf; // 112 * -pi/512
    rom[113] = 32'hbf317fff; // 113 * -pi/512
    rom[114] = 32'hbf33121f; // 114 * -pi/512
    rom[115] = 32'hbf34a43e; // 115 * -pi/512
    rom[116] = 32'hbf36365e; // 116 * -pi/512
    rom[117] = 32'hbf37c87e; // 117 * -pi/512
    rom[118] = 32'hbf395a9e; // 118 * -pi/512
    rom[119] = 32'hbf3aecbd; // 119 * -pi/512
    rom[120] = 32'hbf3c7edd; // 120 * -pi/512
    rom[121] = 32'hbf3e10fd; // 121 * -pi/512
    rom[122] = 32'hbf3fa31c; // 122 * -pi/512
    rom[123] = 32'hbf41353c; // 123 * -pi/512
    rom[124] = 32'hbf42c75c; // 124 * -pi/512
    rom[125] = 32'hbf44597c; // 125 * -pi/512
    rom[126] = 32'hbf45eb9b; // 126 * -pi/512
    rom[127] = 32'hbf477dbb; // 127 * -pi/512
    rom[128] = 32'hbf490fdb; // 128 * -pi/512
    rom[129] = 32'hbf4aa1fa; // 129 * -pi/512
    rom[130] = 32'hbf4c341a; // 130 * -pi/512
    rom[131] = 32'hbf4dc63a; // 131 * -pi/512
    rom[132] = 32'hbf4f5859; // 132 * -pi/512
    rom[133] = 32'hbf50ea79; // 133 * -pi/512
    rom[134] = 32'hbf527c99; // 134 * -pi/512
    rom[135] = 32'hbf540eb9; // 135 * -pi/512
    rom[136] = 32'hbf55a0d8; // 136 * -pi/512
    rom[137] = 32'hbf5732f8; // 137 * -pi/512
    rom[138] = 32'hbf58c518; // 138 * -pi/512
    rom[139] = 32'hbf5a5737; // 139 * -pi/512
    rom[140] = 32'hbf5be957; // 140 * -pi/512
    rom[141] = 32'hbf5d7b77; // 141 * -pi/512
    rom[142] = 32'hbf5f0d97; // 142 * -pi/512
    rom[143] = 32'hbf609fb6; // 143 * -pi/512
    rom[144] = 32'hbf6231d6; // 144 * -pi/512
    rom[145] = 32'hbf63c3f6; // 145 * -pi/512
    rom[146] = 32'hbf655615; // 146 * -pi/512
    rom[147] = 32'hbf66e835; // 147 * -pi/512
    rom[148] = 32'hbf687a55; // 148 * -pi/512
    rom[149] = 32'hbf6a0c75; // 149 * -pi/512
    rom[150] = 32'hbf6b9e94; // 150 * -pi/512
    rom[151] = 32'hbf6d30b4; // 151 * -pi/512
    rom[152] = 32'hbf6ec2d4; // 152 * -pi/512
    rom[153] = 32'hbf7054f3; // 153 * -pi/512
    rom[154] = 32'hbf71e713; // 154 * -pi/512
    rom[155] = 32'hbf737933; // 155 * -pi/512
    rom[156] = 32'hbf750b52; // 156 * -pi/512
    rom[157] = 32'hbf769d72; // 157 * -pi/512
    rom[158] = 32'hbf782f92; // 158 * -pi/512
    rom[159] = 32'hbf79c1b2; // 159 * -pi/512
    rom[160] = 32'hbf7b53d1; // 160 * -pi/512
    rom[161] = 32'hbf7ce5f1; // 161 * -pi/512
    rom[162] = 32'hbf7e7811; // 162 * -pi/512
    rom[163] = 32'hbf800518; // 163 * -pi/512
    rom[164] = 32'hbf80ce28; // 164 * -pi/512
    rom[165] = 32'hbf819738; // 165 * -pi/512
    rom[166] = 32'hbf826048; // 166 * -pi/512
    rom[167] = 32'hbf832958; // 167 * -pi/512
    rom[168] = 32'hbf83f267; // 168 * -pi/512
    rom[169] = 32'hbf84bb77; // 169 * -pi/512
    rom[170] = 32'hbf858487; // 170 * -pi/512
    rom[171] = 32'hbf864d97; // 171 * -pi/512
    rom[172] = 32'hbf8716a7; // 172 * -pi/512
    rom[173] = 32'hbf87dfb7; // 173 * -pi/512
    rom[174] = 32'hbf88a8c7; // 174 * -pi/512
    rom[175] = 32'hbf8971d6; // 175 * -pi/512
    rom[176] = 32'hbf8a3ae6; // 176 * -pi/512
    rom[177] = 32'hbf8b03f6; // 177 * -pi/512
    rom[178] = 32'hbf8bcd06; // 178 * -pi/512
    rom[179] = 32'hbf8c9616; // 179 * -pi/512
    rom[180] = 32'hbf8d5f26; // 180 * -pi/512
    rom[181] = 32'hbf8e2836; // 181 * -pi/512
    rom[182] = 32'hbf8ef145; // 182 * -pi/512
    rom[183] = 32'hbf8fba55; // 183 * -pi/512
    rom[184] = 32'hbf908365; // 184 * -pi/512
    rom[185] = 32'hbf914c75; // 185 * -pi/512
    rom[186] = 32'hbf921585; // 186 * -pi/512
    rom[187] = 32'hbf92de95; // 187 * -pi/512
    rom[188] = 32'hbf93a7a5; // 188 * -pi/512
    rom[189] = 32'hbf9470b4; // 189 * -pi/512
    rom[190] = 32'hbf9539c4; // 190 * -pi/512
    rom[191] = 32'hbf9602d4; // 191 * -pi/512
    rom[192] = 32'hbf96cbe4; // 192 * -pi/512
    rom[193] = 32'hbf9794f4; // 193 * -pi/512
    rom[194] = 32'hbf985e04; // 194 * -pi/512
    rom[195] = 32'hbf992714; // 195 * -pi/512
    rom[196] = 32'hbf99f023; // 196 * -pi/512
    rom[197] = 32'hbf9ab933; // 197 * -pi/512
    rom[198] = 32'hbf9b8243; // 198 * -pi/512
    rom[199] = 32'hbf9c4b53; // 199 * -pi/512
    rom[200] = 32'hbf9d1463; // 200 * -pi/512
    rom[201] = 32'hbf9ddd73; // 201 * -pi/512
    rom[202] = 32'hbf9ea683; // 202 * -pi/512
    rom[203] = 32'hbf9f6f92; // 203 * -pi/512
    rom[204] = 32'hbfa038a2; // 204 * -pi/512
    rom[205] = 32'hbfa101b2; // 205 * -pi/512
    rom[206] = 32'hbfa1cac2; // 206 * -pi/512
    rom[207] = 32'hbfa293d2; // 207 * -pi/512
    rom[208] = 32'hbfa35ce2; // 208 * -pi/512
    rom[209] = 32'hbfa425f1; // 209 * -pi/512
    rom[210] = 32'hbfa4ef01; // 210 * -pi/512
    rom[211] = 32'hbfa5b811; // 211 * -pi/512
    rom[212] = 32'hbfa68121; // 212 * -pi/512
    rom[213] = 32'hbfa74a31; // 213 * -pi/512
    rom[214] = 32'hbfa81341; // 214 * -pi/512
    rom[215] = 32'hbfa8dc51; // 215 * -pi/512
    rom[216] = 32'hbfa9a560; // 216 * -pi/512
    rom[217] = 32'hbfaa6e70; // 217 * -pi/512
    rom[218] = 32'hbfab3780; // 218 * -pi/512
    rom[219] = 32'hbfac0090; // 219 * -pi/512
    rom[220] = 32'hbfacc9a0; // 220 * -pi/512
    rom[221] = 32'hbfad92b0; // 221 * -pi/512
    rom[222] = 32'hbfae5bc0; // 222 * -pi/512
    rom[223] = 32'hbfaf24cf; // 223 * -pi/512
    rom[224] = 32'hbfafeddf; // 224 * -pi/512
    rom[225] = 32'hbfb0b6ef; // 225 * -pi/512
    rom[226] = 32'hbfb17fff; // 226 * -pi/512
    rom[227] = 32'hbfb2490f; // 227 * -pi/512
    rom[228] = 32'hbfb3121f; // 228 * -pi/512
    rom[229] = 32'hbfb3db2f; // 229 * -pi/512
    rom[230] = 32'hbfb4a43e; // 230 * -pi/512
    rom[231] = 32'hbfb56d4e; // 231 * -pi/512
    rom[232] = 32'hbfb6365e; // 232 * -pi/512
    rom[233] = 32'hbfb6ff6e; // 233 * -pi/512
    rom[234] = 32'hbfb7c87e; // 234 * -pi/512
    rom[235] = 32'hbfb8918e; // 235 * -pi/512
    rom[236] = 32'hbfb95a9e; // 236 * -pi/512
    rom[237] = 32'hbfba23ad; // 237 * -pi/512
    rom[238] = 32'hbfbaecbd; // 238 * -pi/512
    rom[239] = 32'hbfbbb5cd; // 239 * -pi/512
    rom[240] = 32'hbfbc7edd; // 240 * -pi/512
    rom[241] = 32'hbfbd47ed; // 241 * -pi/512
    rom[242] = 32'hbfbe10fd; // 242 * -pi/512
    rom[243] = 32'hbfbeda0d; // 243 * -pi/512
    rom[244] = 32'hbfbfa31c; // 244 * -pi/512
    rom[245] = 32'hbfc06c2c; // 245 * -pi/512
    rom[246] = 32'hbfc1353c; // 246 * -pi/512
    rom[247] = 32'hbfc1fe4c; // 247 * -pi/512
    rom[248] = 32'hbfc2c75c; // 248 * -pi/512
    rom[249] = 32'hbfc3906c; // 249 * -pi/512
    rom[250] = 32'hbfc4597c; // 250 * -pi/512
    rom[251] = 32'hbfc5228b; // 251 * -pi/512
    rom[252] = 32'hbfc5eb9b; // 252 * -pi/512
    rom[253] = 32'hbfc6b4ab; // 253 * -pi/512
    rom[254] = 32'hbfc77dbb; // 254 * -pi/512
    rom[255] = 32'hbfc846cb; // 255 * -pi/512
    rom[256] = 32'hbfc90fdb; // 256 * -pi/512
    rom[257] = 32'hbfc9d8ea; // 257 * -pi/512
    rom[258] = 32'hbfcaa1fa; // 258 * -pi/512
    rom[259] = 32'hbfcb6b0a; // 259 * -pi/512
    rom[260] = 32'hbfcc341a; // 260 * -pi/512
    rom[261] = 32'hbfccfd2a; // 261 * -pi/512
    rom[262] = 32'hbfcdc63a; // 262 * -pi/512
    rom[263] = 32'hbfce8f4a; // 263 * -pi/512
    rom[264] = 32'hbfcf5859; // 264 * -pi/512
    rom[265] = 32'hbfd02169; // 265 * -pi/512
    rom[266] = 32'hbfd0ea79; // 266 * -pi/512
    rom[267] = 32'hbfd1b389; // 267 * -pi/512
    rom[268] = 32'hbfd27c99; // 268 * -pi/512
    rom[269] = 32'hbfd345a9; // 269 * -pi/512
    rom[270] = 32'hbfd40eb9; // 270 * -pi/512
    rom[271] = 32'hbfd4d7c8; // 271 * -pi/512
    rom[272] = 32'hbfd5a0d8; // 272 * -pi/512
    rom[273] = 32'hbfd669e8; // 273 * -pi/512
    rom[274] = 32'hbfd732f8; // 274 * -pi/512
    rom[275] = 32'hbfd7fc08; // 275 * -pi/512
    rom[276] = 32'hbfd8c518; // 276 * -pi/512
    rom[277] = 32'hbfd98e28; // 277 * -pi/512
    rom[278] = 32'hbfda5737; // 278 * -pi/512
    rom[279] = 32'hbfdb2047; // 279 * -pi/512
    rom[280] = 32'hbfdbe957; // 280 * -pi/512
    rom[281] = 32'hbfdcb267; // 281 * -pi/512
    rom[282] = 32'hbfdd7b77; // 282 * -pi/512
    rom[283] = 32'hbfde4487; // 283 * -pi/512
    rom[284] = 32'hbfdf0d97; // 284 * -pi/512
    rom[285] = 32'hbfdfd6a6; // 285 * -pi/512
    rom[286] = 32'hbfe09fb6; // 286 * -pi/512
    rom[287] = 32'hbfe168c6; // 287 * -pi/512
    rom[288] = 32'hbfe231d6; // 288 * -pi/512
    rom[289] = 32'hbfe2fae6; // 289 * -pi/512
    rom[290] = 32'hbfe3c3f6; // 290 * -pi/512
    rom[291] = 32'hbfe48d06; // 291 * -pi/512
    rom[292] = 32'hbfe55615; // 292 * -pi/512
    rom[293] = 32'hbfe61f25; // 293 * -pi/512
    rom[294] = 32'hbfe6e835; // 294 * -pi/512
    rom[295] = 32'hbfe7b145; // 295 * -pi/512
    rom[296] = 32'hbfe87a55; // 296 * -pi/512
    rom[297] = 32'hbfe94365; // 297 * -pi/512
    rom[298] = 32'hbfea0c75; // 298 * -pi/512
    rom[299] = 32'hbfead584; // 299 * -pi/512
    rom[300] = 32'hbfeb9e94; // 300 * -pi/512
    rom[301] = 32'hbfec67a4; // 301 * -pi/512
    rom[302] = 32'hbfed30b4; // 302 * -pi/512
    rom[303] = 32'hbfedf9c4; // 303 * -pi/512
    rom[304] = 32'hbfeec2d4; // 304 * -pi/512
    rom[305] = 32'hbfef8be3; // 305 * -pi/512
    rom[306] = 32'hbff054f3; // 306 * -pi/512
    rom[307] = 32'hbff11e03; // 307 * -pi/512
    rom[308] = 32'hbff1e713; // 308 * -pi/512
    rom[309] = 32'hbff2b023; // 309 * -pi/512
    rom[310] = 32'hbff37933; // 310 * -pi/512
    rom[311] = 32'hbff44243; // 311 * -pi/512
    rom[312] = 32'hbff50b52; // 312 * -pi/512
    rom[313] = 32'hbff5d462; // 313 * -pi/512
    rom[314] = 32'hbff69d72; // 314 * -pi/512
    rom[315] = 32'hbff76682; // 315 * -pi/512
    rom[316] = 32'hbff82f92; // 316 * -pi/512
    rom[317] = 32'hbff8f8a2; // 317 * -pi/512
    rom[318] = 32'hbff9c1b2; // 318 * -pi/512
    rom[319] = 32'hbffa8ac1; // 319 * -pi/512
    rom[320] = 32'hbffb53d1; // 320 * -pi/512
    rom[321] = 32'hbffc1ce1; // 321 * -pi/512
    rom[322] = 32'hbffce5f1; // 322 * -pi/512
    rom[323] = 32'hbffdaf01; // 323 * -pi/512
    rom[324] = 32'hbffe7811; // 324 * -pi/512
    rom[325] = 32'hbfff4121; // 325 * -pi/512
    rom[326] = 32'hc0000518; // 326 * -pi/512
    rom[327] = 32'hc00069a0; // 327 * -pi/512
    rom[328] = 32'hc000ce28; // 328 * -pi/512
    rom[329] = 32'hc00132b0; // 329 * -pi/512
    rom[330] = 32'hc0019738; // 330 * -pi/512
    rom[331] = 32'hc001fbc0; // 331 * -pi/512
    rom[332] = 32'hc0026048; // 332 * -pi/512
    rom[333] = 32'hc002c4d0; // 333 * -pi/512
    rom[334] = 32'hc0032958; // 334 * -pi/512
    rom[335] = 32'hc0038de0; // 335 * -pi/512
    rom[336] = 32'hc003f267; // 336 * -pi/512
    rom[337] = 32'hc00456ef; // 337 * -pi/512
    rom[338] = 32'hc004bb77; // 338 * -pi/512
    rom[339] = 32'hc0051fff; // 339 * -pi/512
    rom[340] = 32'hc0058487; // 340 * -pi/512
    rom[341] = 32'hc005e90f; // 341 * -pi/512
    rom[342] = 32'hc0064d97; // 342 * -pi/512
    rom[343] = 32'hc006b21f; // 343 * -pi/512
    rom[344] = 32'hc00716a7; // 344 * -pi/512
    rom[345] = 32'hc0077b2f; // 345 * -pi/512
    rom[346] = 32'hc007dfb7; // 346 * -pi/512
    rom[347] = 32'hc008443f; // 347 * -pi/512
    rom[348] = 32'hc008a8c7; // 348 * -pi/512
    rom[349] = 32'hc0090d4f; // 349 * -pi/512
    rom[350] = 32'hc00971d6; // 350 * -pi/512
    rom[351] = 32'hc009d65e; // 351 * -pi/512
    rom[352] = 32'hc00a3ae6; // 352 * -pi/512
    rom[353] = 32'hc00a9f6e; // 353 * -pi/512
    rom[354] = 32'hc00b03f6; // 354 * -pi/512
    rom[355] = 32'hc00b687e; // 355 * -pi/512
    rom[356] = 32'hc00bcd06; // 356 * -pi/512
    rom[357] = 32'hc00c318e; // 357 * -pi/512
    rom[358] = 32'hc00c9616; // 358 * -pi/512
    rom[359] = 32'hc00cfa9e; // 359 * -pi/512
    rom[360] = 32'hc00d5f26; // 360 * -pi/512
    rom[361] = 32'hc00dc3ae; // 361 * -pi/512
    rom[362] = 32'hc00e2836; // 362 * -pi/512
    rom[363] = 32'hc00e8cbe; // 363 * -pi/512
    rom[364] = 32'hc00ef145; // 364 * -pi/512
    rom[365] = 32'hc00f55cd; // 365 * -pi/512
    rom[366] = 32'hc00fba55; // 366 * -pi/512
    rom[367] = 32'hc0101edd; // 367 * -pi/512
    rom[368] = 32'hc0108365; // 368 * -pi/512
    rom[369] = 32'hc010e7ed; // 369 * -pi/512
    rom[370] = 32'hc0114c75; // 370 * -pi/512
    rom[371] = 32'hc011b0fd; // 371 * -pi/512
    rom[372] = 32'hc0121585; // 372 * -pi/512
    rom[373] = 32'hc0127a0d; // 373 * -pi/512
    rom[374] = 32'hc012de95; // 374 * -pi/512
    rom[375] = 32'hc013431d; // 375 * -pi/512
    rom[376] = 32'hc013a7a5; // 376 * -pi/512
    rom[377] = 32'hc0140c2c; // 377 * -pi/512
    rom[378] = 32'hc01470b4; // 378 * -pi/512
    rom[379] = 32'hc014d53c; // 379 * -pi/512
    rom[380] = 32'hc01539c4; // 380 * -pi/512
    rom[381] = 32'hc0159e4c; // 381 * -pi/512
    rom[382] = 32'hc01602d4; // 382 * -pi/512
    rom[383] = 32'hc016675c; // 383 * -pi/512
    rom[384] = 32'hc016cbe4; // 384 * -pi/512
    rom[385] = 32'hc017306c; // 385 * -pi/512
    rom[386] = 32'hc01794f4; // 386 * -pi/512
    rom[387] = 32'hc017f97c; // 387 * -pi/512
    rom[388] = 32'hc0185e04; // 388 * -pi/512
    rom[389] = 32'hc018c28c; // 389 * -pi/512
    rom[390] = 32'hc0192714; // 390 * -pi/512
    rom[391] = 32'hc0198b9b; // 391 * -pi/512
    rom[392] = 32'hc019f023; // 392 * -pi/512
    rom[393] = 32'hc01a54ab; // 393 * -pi/512
    rom[394] = 32'hc01ab933; // 394 * -pi/512
    rom[395] = 32'hc01b1dbb; // 395 * -pi/512
    rom[396] = 32'hc01b8243; // 396 * -pi/512
    rom[397] = 32'hc01be6cb; // 397 * -pi/512
    rom[398] = 32'hc01c4b53; // 398 * -pi/512
    rom[399] = 32'hc01cafdb; // 399 * -pi/512
    rom[400] = 32'hc01d1463; // 400 * -pi/512
    rom[401] = 32'hc01d78eb; // 401 * -pi/512
    rom[402] = 32'hc01ddd73; // 402 * -pi/512
    rom[403] = 32'hc01e41fb; // 403 * -pi/512
    rom[404] = 32'hc01ea683; // 404 * -pi/512
    rom[405] = 32'hc01f0b0a; // 405 * -pi/512
    rom[406] = 32'hc01f6f92; // 406 * -pi/512
    rom[407] = 32'hc01fd41a; // 407 * -pi/512
    rom[408] = 32'hc02038a2; // 408 * -pi/512
    rom[409] = 32'hc0209d2a; // 409 * -pi/512
    rom[410] = 32'hc02101b2; // 410 * -pi/512
    rom[411] = 32'hc021663a; // 411 * -pi/512
    rom[412] = 32'hc021cac2; // 412 * -pi/512
    rom[413] = 32'hc0222f4a; // 413 * -pi/512
    rom[414] = 32'hc02293d2; // 414 * -pi/512
    rom[415] = 32'hc022f85a; // 415 * -pi/512
    rom[416] = 32'hc0235ce2; // 416 * -pi/512
    rom[417] = 32'hc023c16a; // 417 * -pi/512
    rom[418] = 32'hc02425f1; // 418 * -pi/512
    rom[419] = 32'hc0248a79; // 419 * -pi/512
    rom[420] = 32'hc024ef01; // 420 * -pi/512
    rom[421] = 32'hc0255389; // 421 * -pi/512
    rom[422] = 32'hc025b811; // 422 * -pi/512
    rom[423] = 32'hc0261c99; // 423 * -pi/512
    rom[424] = 32'hc0268121; // 424 * -pi/512
    rom[425] = 32'hc026e5a9; // 425 * -pi/512
    rom[426] = 32'hc0274a31; // 426 * -pi/512
    rom[427] = 32'hc027aeb9; // 427 * -pi/512
    rom[428] = 32'hc0281341; // 428 * -pi/512
    rom[429] = 32'hc02877c9; // 429 * -pi/512
    rom[430] = 32'hc028dc51; // 430 * -pi/512
    rom[431] = 32'hc02940d9; // 431 * -pi/512
    rom[432] = 32'hc029a560; // 432 * -pi/512
    rom[433] = 32'hc02a09e8; // 433 * -pi/512
    rom[434] = 32'hc02a6e70; // 434 * -pi/512
    rom[435] = 32'hc02ad2f8; // 435 * -pi/512
    rom[436] = 32'hc02b3780; // 436 * -pi/512
    rom[437] = 32'hc02b9c08; // 437 * -pi/512
    rom[438] = 32'hc02c0090; // 438 * -pi/512
    rom[439] = 32'hc02c6518; // 439 * -pi/512
    rom[440] = 32'hc02cc9a0; // 440 * -pi/512
    rom[441] = 32'hc02d2e28; // 441 * -pi/512
    rom[442] = 32'hc02d92b0; // 442 * -pi/512
    rom[443] = 32'hc02df738; // 443 * -pi/512
    rom[444] = 32'hc02e5bc0; // 444 * -pi/512
    rom[445] = 32'hc02ec048; // 445 * -pi/512
    rom[446] = 32'hc02f24cf; // 446 * -pi/512
    rom[447] = 32'hc02f8957; // 447 * -pi/512
    rom[448] = 32'hc02feddf; // 448 * -pi/512
    rom[449] = 32'hc0305267; // 449 * -pi/512
    rom[450] = 32'hc030b6ef; // 450 * -pi/512
    rom[451] = 32'hc0311b77; // 451 * -pi/512
    rom[452] = 32'hc0317fff; // 452 * -pi/512
    rom[453] = 32'hc031e487; // 453 * -pi/512
    rom[454] = 32'hc032490f; // 454 * -pi/512
    rom[455] = 32'hc032ad97; // 455 * -pi/512
    rom[456] = 32'hc033121f; // 456 * -pi/512
    rom[457] = 32'hc03376a7; // 457 * -pi/512
    rom[458] = 32'hc033db2f; // 458 * -pi/512
    rom[459] = 32'hc0343fb7; // 459 * -pi/512
    rom[460] = 32'hc034a43e; // 460 * -pi/512
    rom[461] = 32'hc03508c6; // 461 * -pi/512
    rom[462] = 32'hc0356d4e; // 462 * -pi/512
    rom[463] = 32'hc035d1d6; // 463 * -pi/512
    rom[464] = 32'hc036365e; // 464 * -pi/512
    rom[465] = 32'hc0369ae6; // 465 * -pi/512
    rom[466] = 32'hc036ff6e; // 466 * -pi/512
    rom[467] = 32'hc03763f6; // 467 * -pi/512
    rom[468] = 32'hc037c87e; // 468 * -pi/512
    rom[469] = 32'hc0382d06; // 469 * -pi/512
    rom[470] = 32'hc038918e; // 470 * -pi/512
    rom[471] = 32'hc038f616; // 471 * -pi/512
    rom[472] = 32'hc0395a9e; // 472 * -pi/512
    rom[473] = 32'hc039bf25; // 473 * -pi/512
    rom[474] = 32'hc03a23ad; // 474 * -pi/512
    rom[475] = 32'hc03a8835; // 475 * -pi/512
    rom[476] = 32'hc03aecbd; // 476 * -pi/512
    rom[477] = 32'hc03b5145; // 477 * -pi/512
    rom[478] = 32'hc03bb5cd; // 478 * -pi/512
    rom[479] = 32'hc03c1a55; // 479 * -pi/512
    rom[480] = 32'hc03c7edd; // 480 * -pi/512
    rom[481] = 32'hc03ce365; // 481 * -pi/512
    rom[482] = 32'hc03d47ed; // 482 * -pi/512
    rom[483] = 32'hc03dac75; // 483 * -pi/512
    rom[484] = 32'hc03e10fd; // 484 * -pi/512
    rom[485] = 32'hc03e7585; // 485 * -pi/512
    rom[486] = 32'hc03eda0d; // 486 * -pi/512
    rom[487] = 32'hc03f3e94; // 487 * -pi/512
    rom[488] = 32'hc03fa31c; // 488 * -pi/512
    rom[489] = 32'hc04007a4; // 489 * -pi/512
    rom[490] = 32'hc0406c2c; // 490 * -pi/512
    rom[491] = 32'hc040d0b4; // 491 * -pi/512
    rom[492] = 32'hc041353c; // 492 * -pi/512
    rom[493] = 32'hc04199c4; // 493 * -pi/512
    rom[494] = 32'hc041fe4c; // 494 * -pi/512
    rom[495] = 32'hc04262d4; // 495 * -pi/512
    rom[496] = 32'hc042c75c; // 496 * -pi/512
    rom[497] = 32'hc0432be4; // 497 * -pi/512
    rom[498] = 32'hc043906c; // 498 * -pi/512
    rom[499] = 32'hc043f4f4; // 499 * -pi/512
    rom[500] = 32'hc044597c; // 500 * -pi/512
    rom[501] = 32'hc044be03; // 501 * -pi/512
    rom[502] = 32'hc045228b; // 502 * -pi/512
    rom[503] = 32'hc0458713; // 503 * -pi/512
    rom[504] = 32'hc045eb9b; // 504 * -pi/512
    rom[505] = 32'hc0465023; // 505 * -pi/512
    rom[506] = 32'hc046b4ab; // 506 * -pi/512
    rom[507] = 32'hc0471933; // 507 * -pi/512
    rom[508] = 32'hc0477dbb; // 508 * -pi/512
    rom[509] = 32'hc047e243; // 509 * -pi/512
    rom[510] = 32'hc04846cb; // 510 * -pi/512
    rom[511] = 32'hc048ab53; // 511 * -pi/512
end

always @(posedge i_clk) begin
    o_data <= rom[i_addr];
end

endmodule
